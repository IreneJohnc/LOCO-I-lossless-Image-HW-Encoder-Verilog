`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:57:34 12/24/2010 
// Design Name: 
// Module Name:    uarttx 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module uarttx(clk, datain, wrsig, idle, tx); 
input clk;          //UARTʱ�� 
input [7:0] datain; //��Ҫ���͵����� 
input wrsig;        //���������������Ч 
output idle;        //��·״ָ̬ʾ����Ϊ��·æ����Ϊ��·���� 
output tx;          //���������ź� 
reg idle, tx; 
reg send; 
reg wrsigbuf, wrsigrise; 
reg presult; 
reg[7:0] cnt;       //������ 
parameter paritymode = 1'b0; 
//��ⷢ�������Ƿ���Ч 
always @(posedge clk) 
begin 
wrsigbuf <= wrsig; 
wrsigrise <= (~wrsigbuf) & wrsig; 
end 
always @(posedge clk) 
begin 
if (wrsigrise &&  (~idle))  //������������Ч����·Ϊ����ʱ�������µ����ݷ��ͽ��� 
begin 
send <= 1'b1; 
end 
else if(cnt == 8'd176)      //һ֡���Ϸ��ͽ��� 
begin 
send <= 1'b0; 
end 
end 
always @(posedge clk) 
begin 
if(send == 1'b1) 
begin 
case(cnt)       //������ʼλ 
8'd0: 
begin 
tx <= 1'b0; 
idle <= 1'b1; 
cnt <= cnt + 8'd1; 
end 
8'd16: 
begin 
tx <= datain[0];    //�������� 0λ 
presult <= datain[0]^paritymode; 
idle <= 1'b1; 
cnt <= cnt + 8'd1; 
end 
8'd32: 
begin 
tx <= datain[1];    //�������� 1λ 
presult <= datain[1]^presult; 
idle <= 1'b1; 
cnt <= cnt + 8'd1; 
end 
8'd48: 
begin 
tx <= datain[2];    //�������� 2λ 
presult <= datain[2]^presult; idle <= 1'b1; 
cnt <= cnt + 8'd1; 
end 
8'd64: 
begin 
tx <= datain[3];    //�������� 3λ 
presult <= datain[3]^presult; 
idle <= 1'b1; 
cnt <= cnt + 8'd1; 
end 
8'd80: 
begin 
tx <= datain[4];    //�������� 4λ 
presult <= datain[4]^presult; 
idle <= 1'b1; 
cnt <= cnt + 8'd1; 
end 
8'd96: 
begin 
tx <= datain[5];    //�������� 5λ 
presult <= datain[5]^presult; 
idle <= 1'b1; 
cnt <= cnt + 8'd1; 
end 8'd112: 
begin 
tx <= datain[6];    //�������� 6λ 
presult <= datain[6]^presult; 
idle <= 1'b1; 
cnt <= cnt + 8'd1; 
end 
8'd128: 
begin 
tx <= datain[7];    //�������� 7λ 
presult <= datain[7]^presult; 
idle <= 1'b1; 
cnt <= cnt + 8'd1; 
end 
8'd144: 
begin 
tx <= presult;      //������żУ��λ 
presult <= datain[0]^paritymode; 
idle <= 1'b1; 
cnt <= cnt + 8'd1; 
end 
8'd160: 
begin 
tx <= 1'b1;     //����ֹͣλ              idle <= 1'b1; 
cnt <= cnt + 8'd1; 
end 
8'd176: 
begin 
tx <= 1'b1;              
idle <= 1'b0;   //һ֡���Ϸ��ͽ��� 
cnt <= cnt + 8'd1; 
end 
default: 
begin 
cnt <= cnt + 8'd1; 
end 
endcase 
end 
else 
begin 
tx <= 1'b1; 
cnt <= 8'd0; 
idle <= 1'b0; 
end 
end 
endmodule
